module mux8to1 (A, B, C, D, E, F, G, H, sel, Q);

  input A, B, C, D, E, F, G, H;
  input [2:0] sel;
  output Q;

/************ your code **************/


/************************************/

endmodule
