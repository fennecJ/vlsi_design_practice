/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor: Tseng Hsin-Yu (Sylvia) --------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02    ---------------------- //
// ---------------------- priority encoder  ---------------------- // 
/////////////////////////////////////////////////////////////////////

// Module name and I/O port
module encoder(I3,I2,I1,I0,O1,O0);

// Input and output ports declaration
input I3,I2,I1,I0;
output O1,O0;
 
/********* your code ***********/




/******************************/

endmodule
