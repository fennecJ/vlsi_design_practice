module grayscale(color,gray);
  input [23:0] color;
  output [7:0] gray;

/************ your code **************/


/************************************/

endmodule
