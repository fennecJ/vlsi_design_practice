/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor : Michael  ---------------------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02.26 ---------------------- //
// ---------------------- Simple Controller ---------------------- //
/////////////////////////////////////////////////////////////////////

module grayscale(
                 d,
                 q
				);

// ---------------------- input  ---------------------- //
	input [23:0]d;
  
// ---------------------- output ---------------------- //  
	output [7:0]q;

// --------------- below is your design --------------- //
  
endmodule
// ------------------ the end of code ------------------ //
