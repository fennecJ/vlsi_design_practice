/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor : 	KevinLin ----------------------//
// ---------------------- Date : 2019.03    ---------------------- //
// ----------------------      test2        ---------------------- // 
/////////////////////////////////////////////////////////////////////
module test2(out1, 
             out2,
             out3, 
             in1, 
             in2);
            
input  in1, in2;
output out1, out2, out3;

assign out1 = in1 & in2;    //and
assign out2 = in1 | in2;   //or
assign out3 = in1 ^ in2;   //xor

endmodule
