/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor : Michael  ---------------------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02.19 ---------------------- //
// ----------------------  Parametric ReLU  ---------------------- //
/////////////////////////////////////////////////////////////////////


module PRelu(in,out);
				
  // ---------------------- input  ---------------------- //
  input  signed		[`Pixel_DataSize*2:0]	in;
 
  // ---------------------- output ---------------------- //
  output  signed	[`Pixel_DataSize*2:0]	out;

  // ----------------------  reg   ---------------------- //
  reg signed		[`Pixel_DataSize*2:0]	out;
  reg[`Pixel_DataSize*2:0] tmp;
  // ---------------------- Write down Your design below  ---------------------- //
  always @(*) begin
    if(in > 0)begin
    out <= in;
    end
    else begin
    out <= (in>>>6);
    end
  end
  endmodule
